//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:14:54 09/09/2012 
// Design Name: 
// Module Name:    key_codes.vh
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

`define KEY_IDLE  3'd0
`define KEY_UP    3'd1
`define KEY_DOWN  3'd2
`define KEY_LEFT  3'd3
`define KEY_RIGHT 3'd4
`define KEY_FLIP  3'd5
`define KEY_NXT   3'd6
